// Copyright 2016 Tudor Timisescu (verificationgentleman.com)
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//     http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.


class filter_sequence extends amiq_apb_master_base_seq;
  virtual task body();
    amiq_apb_master_simple_seq write_seq;
    `uvm_do_with(write_seq, {
      master_address == 0;
      master_rw == WRITE;
    })
  endtask

  function new(string name = "filter_sequence");
    super.new(name);
  endfunction

  `uvm_object_utils(apb_pipeline_tb::filter_sequence)
endclass
