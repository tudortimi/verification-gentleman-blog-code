// Copyright 2015 Tudor Timisescu (verificationgentleman.com)
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//     http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.


class instruction;
  rand operation_e operation;
  rand register_e op1;
  rand register_e op2;
  rand register_e dest;

  function void print();
    $display("%s %s and %s to %s", operation.name(), op1.name(), op2.name(),
      dest.name());
  endfunction
endclass
