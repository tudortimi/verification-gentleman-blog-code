// Copyright 2014 Tudor Timisescu (verificationgentleman.com)
// 
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
// 
//     http://www.apache.org/licenses/LICENSE-2.0
// 
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.


module top;
  import vgm_uvm_additions_pkg::*;
  
  initial begin
    static vgm_uvm_component comp = new("comp", null);
    static vgm_uvm_monitor mon = new("mon", null);
    
    comp.start_of_simulation_phase(null);
    mon.start_of_simulation_phase(null);
  end
endmodule
