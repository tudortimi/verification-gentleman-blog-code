// Copyright 2014 Tudor Timisescu (verificationgentleman.com)
// 
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
// 
//     http://www.apache.org/licenses/LICENSE-2.0
// 
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.


package example_reg_pkg;
  import uvm_pkg::*;
  `include "uvm_macros.svh"
  
  `include "vgm_rwi0_reg_field.svh"
  
  `include "example_reg_item.svh"
  `include "example_reg_type.svh"
  `include "example_reg_block_type.svh"
  `include "example_reg_test.svh"  
endpackage
