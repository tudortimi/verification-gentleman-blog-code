// Copyright 2016 Tudor Timisescu (verificationgentleman.com)
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//     http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.


package apb_pipeline_tb;
  import uvm_pkg::*;
  `include "uvm_macros.svh"

  import amiq_apb_pkg::*;

  `include "apb_pipeline_tb_scoreboard.svh"
  `include "apb_pipeline_tb_env.svh"
  `include "apb_pipeline_tb_seq_lib.svh"
endpackage
